* D:\OneDrive\Polibuda\KoNaR\1 Linefollower - Projekt\schemat_KiCad\PŁYTKA PRZEDNIA\płytka_przednia.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 14.11.2016 20:12:10

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
T1  Net-_R11-Pad2_ Net-_T1-Pad2_ GND /T1 KTIR0711S		
R11  VCC Net-_R11-Pad2_ 200		
R12  VCC /T1 10K		
T3  Net-_R31-Pad2_ Net-_T3-Pad2_ GND /T3 KTIR0711S		
R31  VCC Net-_R31-Pad2_ 200		
R32  VCC /T3 10k		
T5  Net-_R51-Pad2_ Net-_T5-Pad2_ GND /T5 KTIR0711S		
R51  VCC Net-_R51-Pad2_ 200		
R52  VCC /T5 10k		
T7  Net-_R71-Pad2_ GND GND /T7 KTIR0711S		
R71  VCC Net-_R71-Pad2_ 200		
R72  VCC /T7 10k		
T2  Net-_R21-Pad2_ GND GND /T2 KTIR0711S		
R21  VCC Net-_R21-Pad2_ 200		
R22  VCC /T2 10k		
T4  Net-_R41-Pad2_ Net-_T4-Pad2_ GND /T4 KTIR0711S		
R41  VCC Net-_R41-Pad2_ 200		
R42  VCC /T4 10k		
T6  Net-_R61-Pad2_ GND GND /T6 KTIR0711S		
R61  VCC Net-_R61-Pad2_ 200		
R62  VCC /T6 10k		
T8  Net-_R81-Pad2_ GND GND /T8 KTIR0711S		
R81  VCC Net-_R81-Pad2_ 200		
R82  VCC /T8 10k		
WYJŚCIE_PLYTKA_TYLNIA1  VCC GND /T1 /T2 /T3 /T4 /T5 /T6 /T7 /T8 PIN10		

.end
